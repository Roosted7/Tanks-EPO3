configuration register_logic_synthesised_cfg of register_logic is
   for synthesised
   end for;
end register_logic_synthesised_cfg;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity input_syst_tb is
end input_syst_tb;



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-------------------------------------------------------------------
----------------   tank compare module testbench   ----------------
-------------------------------------------------------------------

-- testbench for module for a subsystem made for epo-3 project at 
--  tu delft
-- project 	: tank game 
-- date		: 25/11/2016
-- subsystem	: pixel generator (aart-peter, niels)
-- author	: aart-peter schipper

-- module computes whether or not to sets of 4 bit x,y coordinates
--  coincide.

-------------------------------------------------------------------

entity tb_tank_comp is
end entity;


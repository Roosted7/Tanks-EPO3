library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of not_gate is
begin
output <= not input;
end behaviour;



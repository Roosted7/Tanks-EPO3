configuration new_pos_vec_behaviour_cfg of new_pos_vec is
   for behaviour
   end for;
end new_pos_vec_behaviour_cfg;



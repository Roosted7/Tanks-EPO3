configuration counter3bit_synthesised_cfg of counter3bit is
   for synthesised
   end for;
end counter3bit_synthesised_cfg;



configuration cfg_beh_pg_pxc of pg_pxc is
   for beh_pg_pxc
   end for;
end cfg_beh_pg_pxc;



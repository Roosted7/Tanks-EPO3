library IEEE;
use IEEE.std_logic_1164.ALL;

entity register1bit is
   port(D  :in    std_logic;
        Q  :out   std_logic;
        clk:in    std_logic;
	reset: in std_logic);
end register1bit;









configuration input_system_synthesised_cfg of input_system is
   for synthesised
      for all: encoder use configuration work.encoder_synthesised_cfg;
      end for;
   end for;
end input_system_synthesised_cfg;



configuration counter3bit_behaviour_cfg of counter3bit is
   for behaviour
   end for;
end counter3bit_behaviour_cfg;



library IEEE;
use IEEE.std_logic_1164.ALL;
use ieee.numeric_std.all;

entity input_fsm_tb is
end input_fsm_tb;






configuration new_top_extracted_cfg of new_top is
   for extracted
   end for;
end new_top_extracted_cfg;



configuration cfg_syn_pg_prg of pg_prg is
   for synthesised
   end for;
end cfg_syn_pg_prg;



configuration tank_pos_reg_synthesised_cfg of tank_pos_reg is
   for synthesised
   end for;
end tank_pos_reg_synthesised_cfg;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity test_logic_2 is
   port(c_5 :in    std_logic;
        c_4 :in    std_logic;
        c_3 :in    std_logic;
        c_2 :in    std_logic;
        c_1 :in    std_logic;
        c_0 :in    std_logic;
        t_e :in    std_logic_vector(2 downto 0);
        pass:out   std_logic);
end test_logic_2;



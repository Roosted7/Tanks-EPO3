configuration register_logic_extracted_cfg of register_logic is
   for extracted
   end for;
end register_logic_extracted_cfg;



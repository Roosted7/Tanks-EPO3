configuration encoder_tb_behaviour_cyn_cfg of encoder_tb is
   for behaviour
      for all: encoder use configuration work.encoder_synthesised_cfg;
      end for;
   end for;
end encoder_tb_behaviour_cyn_cfg;



configuration cfg_pix_comp of pix_comp is
   for beh_pix_comp
   end for;
end cfg_pix_comp;



library IEEE;
use IEEE.std_logic_1164.ALL;

architecture beh_tank_hr of tank_hit_reg is
begin

process (clk, reset)
	if (rising_edge(clk)) then
		

end beh_tank_hr;



configuration combiblok_coord_tb_behaviour_cfg of combiblok_coord_tb is
   for behaviour
      for all: combiblok_coord use configuration work.combiblok_coord_behaviour_cfg;
      end for;
   end for;
end combiblok_coord_tb_behaviour_cfg;



configuration tank_pos_reg_extracted_cfg of tank_pos_reg is
   for extracted
   end for;
end tank_pos_reg_extracted_cfg;



configuration register1bit_synthesised_cfg of register1bit is
   for synthesised
   end for;
end register1bit_synthesised_cfg;



configuration new_pos_vec_extracted_cfg of new_pos_vec is
   for extracted
   end for;
end new_pos_vec_extracted_cfg;



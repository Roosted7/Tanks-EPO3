library IEEE;
use IEEE.std_logic_1164.ALL;

entity new_pos_vec_tb is
end new_pos_vec_tb;



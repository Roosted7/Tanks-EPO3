configuration encoder_tb_behaviour_cfg of encoder_tb is
   for behaviour
      for all: encoder use configuration work.encoder_behaviour_cfg;
      end for;
   end for;
end encoder_tb_behaviour_cfg;



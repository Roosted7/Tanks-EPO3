configuration new_coord_tb_behaviour_cfg of new_coord_tb is
   for behaviour
      for all: new_coord use configuration work.new_coord_structural_cfg;
      end for;
   end for;
end new_coord_tb_behaviour_cfg;



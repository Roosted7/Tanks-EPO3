configuration input_system_extracted_cfg of input_system is
   for extracted
   end for;
end input_system_extracted_cfg;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity counter3bit is
    Port ( CLK : in  STD_LOGIC;
           Count : out  STD_LOGIC_VECTOR (2 downto 0));
end counter3bit;





configuration tf_rise_behaviour_cfg of tf_rise is
   for behaviour
   end for;
end tf_rise_behaviour_cfg;



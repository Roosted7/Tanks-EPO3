library IEEE;
use IEEE.std_logic_1164.ALL;

entity input_fsm_tb is
end input_fsm_tb;



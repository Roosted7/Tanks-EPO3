configuration tb_beh_top_1 of tb_pg_top is
   for beh_top
      for all: pg_top use configuration work.pg_player_1;
      end for;
   end for;
end tb_beh_top_1;



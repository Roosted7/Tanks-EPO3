configuration cfg_syn_pg_hrg of pg_hrg is
   for synthesised
   end for;
end cfg_syn_pg_hrg;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity tf_rise is
   port(tf_in  :in    std_logic;
	reset  :in	   std_logic;
	clk    :in    std_logic;
        tf_rise:out   std_logic);
end tf_rise;






configuration cfg_ext_pg_tkc of pg_tkc is
   for extracted
   end for;
end cfg_ext_pg_tkc;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity newposition_tb is
end newposition_tb;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity audio is
   port(clk_30     :in    std_logic;
        clk_30k    :in    std_logic;
        reset		   :in    std_logic;
        music      :out   std_logic);
end audio;






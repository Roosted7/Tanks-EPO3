library IEEE;
use IEEE.std_logic_1164.ALL;

entity input_reg_tb is
end input_reg_tb;



configuration register_logic_behaviour_cfg of register_logic is
   for behaviour
   end for;
end register_logic_behaviour_cfg;



configuration cfg_ext_pg_hrg of pg_hrg is
   for extracted
   end for;
end cfg_ext_pg_hrg;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity test_clear is
   port(input :in    std_logic;
	test_enable: in std_logic;
        clk   :in    std_logic;
        reset :in    std_logic;
        output:out   std_logic);
end test_clear;






library IEEE;
use IEEE.std_logic_1164.ALL;

entity s is
   port(inp :in    std_logic_vector(2 downto 0);
        outp:out   std_logic);
end s;












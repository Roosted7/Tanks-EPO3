library IEEE;
use IEEE.std_logic_1164.ALL;

entity tl_pg_tank is
end tl_pg_tank;



configuration calculated_new_pos_tb_behaviour_cfg of calculated_new_pos_tb is
   for behaviour
      for all: calculated_new_pos use configuration work.calculated_new_pos_structural_cfg;
      end for;
   end for;
end calculated_new_pos_tb_behaviour_cfg;



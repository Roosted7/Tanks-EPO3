library IEEE;
use IEEE.std_logic_1164.ALL;

entity pulse is
   port(clk    :in    std_logic;
        bulletd:in    std_logic;
        bulletc:in    std_logic;
        pulse  :out   std_logic);
end pulse;






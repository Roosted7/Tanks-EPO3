configuration input_fsm_behaviour_cfg of input_fsm is
   for behaviour
   end for;
end input_fsm_behaviour_cfg;



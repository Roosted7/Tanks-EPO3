library IEEE;
use IEEE.std_logic_1164.ALL;

entity tb_pg_pxc is
end tb_pg_pxc;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity reg_tb is
end reg_tb;



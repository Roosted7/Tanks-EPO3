library IEEE;
use IEEE.std_logic_1164.ALL;

entity adder_5bits_tb is
end adder_5bits_tb;



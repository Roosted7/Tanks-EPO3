library IEEE;
use IEEE.std_logic_1164.ALL;

entity combiblok_coord_tb is
end combiblok_coord_tb;



configuration combiblok_coord_synthesised_cfg of combiblok_coord is
   for synthesised
   end for;
end combiblok_coord_synthesised_cfg;



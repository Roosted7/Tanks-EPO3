configuration cfg_pg_tank of tl_pg_tank is
   for beh_pg_tank
   end for;
end cfg_pg_tank;



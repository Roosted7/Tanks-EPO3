configuration mux_8bits_synthesised_cfg of mux_8bits is
   for synthesised
   end for;
end mux_8bits_synthesised_cfg;



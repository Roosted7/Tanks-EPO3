library ieee;
use ieee.std_logic_1164.all;

architecture beh_tank_pg of tank_pg is
	-- Memory for the middle pixel of the tank and its orientation.
	-- Uses rising edge of the screen-refresh
	
	component tank_pos_reg is
		port(
			tank_x_in 	: in std_logic_vector(3 downto 0);
			tank_x_out : out std_logic_vector(3 downto 0);
			tank_y_in  : in std_logic_vector(3 downto 0);
			tank_y_out : out std_logic_vector(3 downto 0);
			tank_or_in : in std_logic_vector(1 downto 0);
			tank_or_out: out std_logic_vector(1 downto 0);
			update_pos : in std_logic
		);
	end component;
		
	-- Memory for the hit-status of the tank. Determines if the tank is dead		, or alive.
	-- Uses rising edge of the clock

	component tank_hit_reg is
		port(
			hit_in : in std_logic;
			hit_out : out std_logic;
			clk : in std_logic
		);
	end component;

	-- Generates the tank based off of its middle pixel and the orientation.
	
	component tank_pix is
		port(
			x_in 	     :in    std_logic_vector(3 downto 0);
			y_in 	     :in    std_logic_vector(3 downto 0);
			theta	     :in    std_logic_vector(1 downto 0);
			x_head  	    :out   std_logic_vector(3 downto 0);
			y_head       :out   std_logic_vector(3 downto 0);
			x_body       :out   std_logic_vector(3 downto 0);
			y_body       :out   std_logic_vector(3 downto 0);
			x_left_leg   :out   std_logic_vector(3 downto 0);
			y_left_leg   :out   std_logic_vector(3 downto 0);
			x_right_leg  :out   std_logic_vector(3 downto 0);
			y_right_leg  :out   std_logic_vector(3 downto 0);
			x_left_foot  :out   std_logic_vector(3 downto 0);
			y_left_foot  :out   std_logic_vector(3 downto 0);
			x_right_foot :out   std_logic_vector(3 downto 0);
			y_right_foot :out   std_logic_vector(3 downto 0)
		);
	end component;

	-- Compares the current screen pixel (x,y), with the individual componen		ts of the tank
	-- which are generated by tank_pix	

	component tank_comp is
		port(
			screen_x_in  :in   std_logic_vector(3 downto 0);
			screen_y_in	 :in   std_logic_vector(3 downto 0);
			x_head       :in   std_logic_vector(3 downto 0);
			y_head       :in   std_logic_vector(3 downto 0);
			x_body       :in   std_logic_vector(3 downto 0);
			y_body       :in   std_logic_vector(3 downto 0);
			x_left_leg   :in   std_logic_vector(3 downto 0);
			y_left_leg   :in   std_logic_vector(3 downto 0);
			x_right_leg  :in   std_logic_vector(3 downto 0);
			y_right_leg  :in   std_logic_vector(3 downto 0);
			x_left_foot  :in   std_logic_vector(3 downto 0);
			y_left_foot  :in   std_logic_vector(3 downto 0);
			x_right_foot :in   std_logic_vector(3 downto 0);
			y_right_foot :in   std_logic_vector(3 downto 0);
			draw_out     :out  std_logic
		);
	end component;

	-- Intermediate signals:
	signal tank_x_q, tank_y_q : std_logic_vector(3 downto 0);
	signal tank_or_q : std_logic_vector(1 downto 0);

	signal x_head, y_head,
	x_body, y_body,
   	x_left_leg, y_left_leg,
   	x_right_leg, y_right_leg,
   	x_left_foot, y_left_foot,
   	x_right_foot, y_right_foot	: std_logic_vector(3 downto 0);

	signal draw_out : std_logic;
	signal hit_out_q : std_logic;
begin

c00: tank_pos_reg port map (
							tank_x_in => tank_x_in,
							tank_x_out => tank_x_q,
							tank_y_in => tank_y_in,
							tank_y_out => tank_y_q,
							tank_or_in => tank_or_in,
							tank_or_out => tank_or_q,
							update_pos => update_pos
						   );
c01: tank_hit_reg port map (
							hit_in => hit_in,
							hit_out => hit_out_q,
							clk => clk
						   );
c02: tank_pix port map (
						x_in => screen_x_in,
						y_in => screen_y_in,
						theta => tank_or_q,
						x_head => x_head, 
						y_head => y_head, 
						x_body => x_body, 
						y_body => y_body, 
						x_left_leg => x_left_leg, 
						y_left_leg => y_left_leg, 
						x_right_leg => x_right_leg, 
						y_right_leg => y_right_leg, 
						x_left_foot => x_left_foot, 
						y_left_foot => y_left_foot, 
						x_right_foot => x_right_foot, 
						y_right_foot => y_right_foot 
					   );
c03: tank_comp port map (
						screen_x_in => screen_x_in,
						screen_y_in => screen_y_in,
						x_head => x_head, 
						y_head => y_head, 
						x_body => x_body, 
						y_body => y_body, 
						x_left_leg => x_left_leg, 
						y_left_leg => y_left_leg, 
						x_right_leg => x_right_leg, 
						y_right_leg => y_right_leg, 
						x_left_foot => x_left_foot, 
						y_left_foot => y_left_foot, 
						x_right_foot => x_right_foot, 
						y_right_foot => y_right_foot,
						draw_out => draw_out
						);

s00: tank_x_out <= tank_x_q;
s01: tank_y_out<= tank_y_q;
s02: tank_or_out<= tank_or_q;
s03: draw <= draw_out and not hit_out_q;
s04: hit_out <= hit_out_q;

end beh_tank_pg;



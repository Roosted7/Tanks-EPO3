configuration tank_pos_top_level_extracted_cfg of tank_pos_top_level is
   for extracted
   end for;
end tank_pos_top_level_extracted_cfg;



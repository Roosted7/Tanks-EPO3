configuration new_pos_vec_tb_behaviour_cfg of new_pos_vec_tb is
   for behaviour
      for all: new_pos_vec use configuration work.new_pos_vec_behaviour_cfg;
      end for;
   end for;
end new_pos_vec_tb_behaviour_cfg;



configuration tb_beh_pxg of tb_pg_pxg is
   for beh_pxg
      for all: pg_pxg use configuration work.cfg_beh_pg_pxg;
      end for;
   end for;
end tb_beh_pxg;



configuration input_fsm_extracted_cfg of input_fsm is
   for extracted
   end for;
end input_fsm_extracted_cfg;



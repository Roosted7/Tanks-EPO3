configuration input_system_behaviour_cfg of input_system is
   for behaviour
      for all: encoder use configuration work.encoder_behaviour_cfg;
      end for;
   end for;
end input_system_behaviour_cfg;



configuration cfg_ext_pg_fsm of pg_fsm is
   for extracted
   end for;
end cfg_ext_pg_fsm;



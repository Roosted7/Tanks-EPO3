configuration c_tank_hit_reg of tank_hit_reg is
   for b_tank_hit_reg
   end for;
end c_tank_hit_reg;



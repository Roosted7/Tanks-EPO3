configuration player_2 of pg_prg is
   for beh_pg_prg_2
   end for;
end player_2;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity gen_bullet is
   port(fire_b1: in    std_logic_vector(2 downto 0);
        tank_b1	:	in	std_logic_vector(10 downto 0);
	gen_b1	: out	std_logic_vector(10 downto 0)); 
end gen_bullet;









library IEEE;
use IEEE.std_logic_1164.ALL;

entity tb_timing is
end tb_timing;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity pass_gate is
   port(input :in    std_logic;
        output:out   std_logic);
end pass_gate;



configuration tank_hit_reg_extracted_cfg of tank_hit_reg is
   for extracted
   end for;
end tank_hit_reg_extracted_cfg;



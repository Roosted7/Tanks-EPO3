configuration cfg_ext_pg_pxc of pg_pxc is
   for extracted
   end for;
end cfg_ext_pg_pxc;



configuration mux_8bits_behaviour_cfg of mux_8bits is
   for behaviour
   end for;
end mux_8bits_behaviour_cfg;



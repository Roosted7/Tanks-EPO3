configuration adder_5bits_extracted_cfg of adder_5bits is
   for extracted
   end for;
end adder_5bits_extracted_cfg;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity toplvl_tb is
end toplvl_tb;



configuration fa_5_bit_synthesised_cfg of fa_5_bit is
   for synthesised
   end for;
end fa_5_bit_synthesised_cfg;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity new_coord_tb is
end new_coord_tb;



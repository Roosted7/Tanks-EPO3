configuration mux_1bits_behaviour_cfg of mux_1bits is
   for behaviour
   end for;
end mux_1bits_behaviour_cfg;



configuration new_pos_vec_synthesised_cfg of new_pos_vec is
   for synthesised
   end for;
end new_pos_vec_synthesised_cfg;



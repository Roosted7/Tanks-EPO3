configuration tf_rise_synthesised_cfg of tf_rise is
   for synthesised
   end for;
end tf_rise_synthesised_cfg;



configuration fa_5_bit_behavioural_cfg of fa_5_bit is
   for behavioural
   end for;
end fa_5_bit_behavioural_cfg;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity reg_logic_tb is
end reg_logic_tb;



configuration tank_hit_reg_synthesised_cfg of tank_hit_reg is
   for synthesised
   end for;
end tank_hit_reg_synthesised_cfg;



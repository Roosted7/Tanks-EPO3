configuration cfg_ext_pg_pxg of pg_pxg is
   for extracted
   end for;
end cfg_ext_pg_pxg;



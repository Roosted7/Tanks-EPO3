configuration cfg_ext_pg_top of pg_top is
   for extracted
   end for;
end cfg_ext_pg_top;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity s_inv is
   port(inp :in    std_logic;
        outp:out   std_logic_vector(2 downto 0));
end s_inv;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity fa_5_bit is
   port(a    :in    std_logic_vector(3 downto 0);
		b	: in std_logic_vector(3 downto 0);
		c 	: out std_logic_vector(4 downto 0)
	);
end fa_5_bit;









configuration tb_beh_tkc of tb_pg_tkc is
   for beh_tkc
      for all: pg_tkc use configuration work.cfg_str_pg_tkc;
      end for;
   end for;
end tb_beh_tkc;



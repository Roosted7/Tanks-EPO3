library IEEE;
use IEEE.std_logic_1164.ALL;

entity del_bullet_tb is
end del_bullet_tb;



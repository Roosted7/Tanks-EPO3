library IEEE;
use IEEE.std_logic_1164.ALL;


-------------------------------------------------------------------
---------------   pixel compare module testbench   ----------------
-------------------------------------------------------------------

-- testbench for module for  a subsystem made for epo-3 project at 
--  tu delft
-- project 	: tank game 
-- date		: 25/11/2016
-- subsystem	: pixel generator (aart-peter, niels)
-- author	: aart-peter schipper

-- module computes whether or not to sets of 4 bit x,y coordinates
--  coincide.

-------------------------------------------------------------------

entity tb_pix_comp is
end tb_pix_comp;



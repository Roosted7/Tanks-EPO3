configuration cfg_tb_pix_c of tb_pix_comp is
   for beh_tb_pix_c
      for all: pix_comp use configuration work.cfg_pix_comp;
      end for;
   end for;
end cfg_tb_pix_c;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity bullet_col_tb is
end bullet_col_tb;



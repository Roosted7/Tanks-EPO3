library IEEE;
use IEEE.std_logic_1164.ALL;

entity test_logic_1 is
   port(c_5:in    std_logic;
        c_4:in    std_logic;
        c_3:in    std_logic;
        c_2:in    std_logic;
        c_1:in    std_logic;
        c_0:in    std_logic;
        p_l:out   std_logic;
        p_r:out   std_logic;
        p_u:out   std_logic;
        p_d:out   std_logic;
        p_f:out   std_logic;
        tf :out   std_logic);
end test_logic_1;









configuration cfg_beh_pg_pxg of pg_pxg is
   for beh_pg_pxg
   end for;
end cfg_beh_pg_pxg;



configuration c_tank_pos_reg of tank_pos_reg is
   for b_tank_pos_reg
   end for;
end c_tank_pos_reg;



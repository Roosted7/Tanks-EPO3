configuration cfg_syn_pg_fsm of pg_fsm is
   for synthesised
   end for;
end cfg_syn_pg_fsm;



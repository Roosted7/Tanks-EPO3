library IEEE;
use IEEE.std_logic_1164.ALL;

entity tff is
   port(reset:in	   std_logic;
	t    :in    std_logic;
        q    :out   std_logic);
end entity tff;












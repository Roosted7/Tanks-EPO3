configuration tankwalls_synthesised_cfg of tankwalls is
   for synthesised
   end for;
end tankwalls_synthesised_cfg;



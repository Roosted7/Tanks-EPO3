configuration input_fsm_synthesised_cfg of input_fsm is
   for synthesised
   end for;
end input_fsm_synthesised_cfg;



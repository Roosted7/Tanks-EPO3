configuration mux_2bits_synthesised_cfg of mux_2bits is
   for synthesised
   end for;
end mux_2bits_synthesised_cfg;



configuration encoder_behaviour_cfg of encoder is
   for behaviour
   end for;
end encoder_behaviour_cfg;



configuration cfg_syn_pg_pxc of pg_pxc is
   for synthesised
   end for;
end cfg_syn_pg_pxc;



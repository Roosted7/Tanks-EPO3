library IEEE;
use IEEE.std_logic_1164.ALL;

entity mux_1bits is
   port(new_1  :out   std_logic;
        old_1  :in    std_logic;
        old_2  :in    std_logic;
        control:in    std_logic);
end mux_1bits;



















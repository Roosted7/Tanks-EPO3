configuration encoder_synthesised_cfg of encoder is
   for synthesised
   end for;
end encoder_synthesised_cfg;



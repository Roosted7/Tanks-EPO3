configuration combiblok_coord_behaviour_cfg of combiblok_coord is
   for behaviour
   end for;
end combiblok_coord_behaviour_cfg;



library IEEE;
use IEEE.std_logic_1164.ALL;

architecture beh_pg_tank of tl_pg_tank is
begin
end beh_pg_tank;



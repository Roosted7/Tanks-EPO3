configuration tf_rise_extracted_cfg of tf_rise is
   for extracted
   end for;
end tf_rise_extracted_cfg;



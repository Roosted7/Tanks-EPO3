library IEEE;
use IEEE.std_logic_1164.ALL;
use ieee.numeric_std.all;

entity input_syst_tb is
end input_syst_tb;






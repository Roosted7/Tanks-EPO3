configuration input_register_behaviour_cfg of input_register is
   for behaviour
   end for;
end input_register_behaviour_cfg;



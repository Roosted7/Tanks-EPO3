configuration cfg_beh_pg_hrg of pg_hrg is
   for beh_pg_hrg
   end for;
end cfg_beh_pg_hrg;



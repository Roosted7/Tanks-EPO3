configuration tb_beh_pxc of tb_pg_pxc is
   for beh_pxc
      for all: pg_pxc use configuration work.cfg_beh_pg_pxc;
      end for;
   end for;
end tb_beh_pxc;



configuration cfg_tank_pix of tank_pix is
   for beh_tank_pix
   end for;
end cfg_tank_pix;



configuration adder_5bits_synthesised_cfg of adder_5bits is
   for synthesised
   end for;
end adder_5bits_synthesised_cfg;



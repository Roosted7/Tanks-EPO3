configuration tb_beh_top_2 of tb_pg_top is
   for beh_top
      for all: pg_top use configuration work.pg_player_2;
      end for;
   end for;
end tb_beh_top_2;



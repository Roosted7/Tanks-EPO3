configuration tankwalls_behaviour_cfg of tankwalls is
   for behaviour
   end for;
end tankwalls_behaviour_cfg;



configuration adder_5bits_behaviour_cfg of adder_5bits is
   for behaviour
   end for;
end adder_5bits_behaviour_cfg;



configuration cfg_ext_pg_prg of pg_prg is
   for extracted
   end for;
end cfg_ext_pg_prg;



configuration player_1 of pg_prg is
   for beh_pg_prg_1
   end for;
end player_1;



configuration newposition_behaviour_cfg of newposition is
   for behaviour
   end for;
end newposition_behaviour_cfg;



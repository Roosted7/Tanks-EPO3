configuration register1bit_behaviour_cfg of register1bit is
   for behaviour
   end for;
end register1bit_behaviour_cfg;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity tankwalls is
   port(coord :in    std_logic_vector(7 downto 0);
        result:out   std_logic);
end tankwalls;



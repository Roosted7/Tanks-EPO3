configuration cfg_beh_pg_fsm of pg_fsm is
   for beh_pg_fsm
   end for;
end cfg_beh_pg_fsm;



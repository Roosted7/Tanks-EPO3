configuration cfg_syn_pg_pxg of pg_pxg is
   for synthesised
   end for;
end cfg_syn_pg_pxg;



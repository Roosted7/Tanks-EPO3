configuration input_register_extracted_cfg of input_register is
   for extracted
   end for;
end input_register_extracted_cfg;



configuration adder_5bits_tb_behaviour_cfg of adder_5bits_tb is
   for behaviour
      for all: adder_5bits use configuration work.adder_5bits_behaviour_cfg;
      end for;
   end for;
end adder_5bits_tb_behaviour_cfg;



library IEEE;
use IEEE.std_logic_1164.ALL;

entity calculated_new_pos_tb is
end calculated_new_pos_tb;



configuration mux_1bits_synthesised_cfg of mux_1bits is
   for synthesised
   end for;
end mux_1bits_synthesised_cfg;



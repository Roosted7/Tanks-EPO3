library IEEE;
use IEEE.std_logic_1164.ALL;

entity tf_rise_tb is
end tf_rise_tb;



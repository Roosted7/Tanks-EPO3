library IEEE;
use IEEE.std_logic_1164.ALL;

entity input_count_tb is
end input_count_tb;



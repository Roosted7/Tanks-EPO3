configuration cfg_tank_pg of tank_pg is
   for beh_tank_pg
   end for;
end cfg_tank_pg;



configuration input_register_synthesised_cfg of input_register is
   for synthesised
   end for;
end input_register_synthesised_cfg;



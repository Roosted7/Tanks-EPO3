library IEEE;
use IEEE.std_logic_1164.ALL;

architecture beh_pg_ prg1 of pg_prg is
begin
end beh_pg_ prg1;


